`timescale 1ns / 1ns
module SMP (input PIN,output pout);
// pin   PIN is      MGTREFCLK0P_115 bank 115 bus_bmb7_J4[0]         H6
//assign PIN=0;
assign pout=PIN;
endmodule
