`timescale 1ns / 1ns

module BUFIO (
	output O,
	input I
);
	buf b(O, I);
endmodule
