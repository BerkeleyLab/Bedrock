module BUFR (input CE, output O, input I);
	buf b(O, I);
endmodule
