module OBUF (output O, input I);
	buf b(O, I);
endmodule
