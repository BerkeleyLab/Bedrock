// ------------------------------------
// COMMS_PACK.VH
// Helper constants for comms_top.v
// ------------------------------------

localparam LBUS_ADDR_WIDTH = 24;
localparam LBUS_DATA_WIDTH = 32;

localparam GTX_ETH_WIDTH   = 20;
localparam GTX_CC_WIDTH    = 16;


