module IDELAYCTRL (
    input  RST,
    input  REFCLK,
    output RDY
);
assign RDY = 1'b1;
endmodule
