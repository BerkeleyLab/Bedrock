// Hand-generated
// Somewhat compatible with machine-generated freq.vh from FERMI builds
`define COHERENT_DEN (7)
`define RF_NUM (1)
// floor(32768*0.5*sec(2*pi*1/7/2)+0.5)
`define AFTERBURNER_COEFF (18185)
// needed by interpon.v to even pass syntax checks
`define CIC_CNTW (6)
`define CIC_PERIOD (14)
`define CIC_MULT 16'd0
