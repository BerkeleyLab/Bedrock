module BUFH (output O, input I);
	buf b(O, I);
endmodule
