`timescale 1ns / 1ns

module BUFG (
	output O,
	input I
);
	buf b(O, I);
endmodule
