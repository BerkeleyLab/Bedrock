module IBUF (output O, input I);
	buf b(O, I);
endmodule
