// !!! Placeholder only !!!

module MMCME4_ADV #(
    parameter BANDWIDTH = "OPTIMIZED",
    parameter real CLKFBOUT_MULT_F = 5.0,
    parameter real CLKFBOUT_PHASE = 0.0,
    parameter CLKFBOUT_USE_FINE_PS = "FALSE",
    parameter real CLKIN1_PERIOD = 0.0,
    parameter real CLKIN2_PERIOD = 0.0,
    parameter real CLKOUT0_DIVIDE_F = 1.0,
    parameter real CLKOUT0_DUTY_CYCLE = 0.5,
    parameter real CLKOUT0_PHASE = 0.0,
    parameter CLKOUT0_USE_FINE_PS = "FALSE",
    parameter integer CLKOUT1_DIVIDE = 1,
    parameter real CLKOUT1_DUTY_CYCLE = 0.5,
    parameter real CLKOUT1_PHASE = 0.0,
    parameter CLKOUT1_USE_FINE_PS = "FALSE",
    parameter integer CLKOUT2_DIVIDE = 1,
    parameter real CLKOUT2_DUTY_CYCLE = 0.5,
    parameter real CLKOUT2_PHASE = 0.0,
    parameter CLKOUT2_USE_FINE_PS = "FALSE",
    parameter integer CLKOUT3_DIVIDE = 1,
    parameter real CLKOUT3_DUTY_CYCLE = 0.5,
    parameter real CLKOUT3_PHASE = 0.0,
    parameter CLKOUT3_USE_FINE_PS = "FALSE",
    parameter CLKOUT4_CASCADE = "FALSE",
    parameter integer CLKOUT4_DIVIDE = 1,
    parameter real CLKOUT4_DUTY_CYCLE = 0.5,
    parameter real CLKOUT4_PHASE = 0.0,
    parameter CLKOUT4_USE_FINE_PS = "FALSE",
    parameter integer CLKOUT5_DIVIDE = 1,
    parameter real CLKOUT5_DUTY_CYCLE = 0.5,
    parameter real CLKOUT5_PHASE = 0.0,
    parameter CLKOUT5_USE_FINE_PS = "FALSE",
    parameter integer CLKOUT6_DIVIDE = 1,
    parameter real CLKOUT6_DUTY_CYCLE = 0.5,
    parameter real CLKOUT6_PHASE = 0.0,
    parameter CLKOUT6_USE_FINE_PS = "FALSE",
    parameter COMPENSATION = "AUTO",
    parameter integer DIVCLK_DIVIDE = 1,
    parameter IS_CLKFBIN_INVERTED = 1'b0,
    parameter IS_CLKIN1_INVERTED = 1'b0,
    parameter IS_CLKIN2_INVERTED = 1'b0,
    parameter IS_CLKINSEL_INVERTED = 1'b0,
    parameter IS_PSEN_INVERTED = 1'b0,
    parameter IS_PSINCDEC_INVERTED = 1'b0,
    parameter IS_PWRDWN_INVERTED = 1'b0,
    parameter IS_RST_INVERTED = 1'b0,
    parameter real REF_JITTER1 = 0.0,
    parameter real REF_JITTER2 = 0.0,
    parameter SS_EN = "FALSE",
    parameter SS_MODE = "CENTER_HIGH",
    parameter integer SS_MOD_PERIOD = 10000,
    parameter STARTUP_WAIT = "FALSE"
)(
    output  CLKFBOUT,
    output  CLKFBOUTB,
    output  CLKOUT0,
    output  CLKOUT0B,
    output  CLKOUT1,
    output  CLKOUT1B,
    output  CLKOUT2,
    output  CLKOUT2B,
    output  CLKOUT3,
    output  CLKOUT3B,
    output  CLKOUT4,
    output  CLKOUT5,
    output  CLKOUT6,
    output  LOCKED,
    input   CLKFBIN,
    input   CLKIN1,
    input   CLKIN2,
    input   CLKINSEL,
    input   PWRDWN,
    input   RST,
    input   DADDR,
    input   DCLK,
    input   DEN,
    input   DI,
    input   DO,
    input   DRDY,
    input   DWE,
    output  CDDCDONE,
    input   CDDCREQ,
    input   PSCLK,
    input   PSEN,
    input   PSINCDEC,
    output  PSDONE,
    output  CLKINSTOPPED,
    output  CLKFBSTOPPED
);

assign CLKOUT0 = CLKIN1;
assign CLKOUT1 = CLKIN1;

endmodule // MMCME2_BASE
