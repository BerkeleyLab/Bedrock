// ------------------------------------
// chitchat_pack.vh
// Shared constants for Chitchat IP
// ------------------------------------

localparam CC_GATEWARE_TYPE = 0;
localparam CC_PROTOCOL_CAT = 6;
localparam CC_PROTOCOL_VER = 1;
localparam CC_K28_5 = 8'b10111100;
