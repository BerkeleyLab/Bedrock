module BUFG (output O, input I);
	buf b(O, I);
endmodule
