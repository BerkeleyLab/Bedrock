module BUFIO (output O, input I);
	buf b(O, I);
endmodule
