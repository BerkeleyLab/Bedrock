module NXP_74AVC4T245 (
	output DIR,
	input dirin
);
assign DIR=dirin;
endmodule
