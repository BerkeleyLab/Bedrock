// ------------------------------------
// COMMS_PACK.VH
// Helper constants for comms_top.v
// ------------------------------------

localparam GTX_ETH_WIDTH   = 20;
localparam GTX_CC_WIDTH    = 16;
