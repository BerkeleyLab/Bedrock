// Software-accessible features for support of digitizer board
// Please keep this as simulatable and portable Verilog!
// Purposefully does not include:
//   adc_test
//   iq_trace
//   slow readout chain (and therefore not adc minmax?)
module digitizer_config(

	// local bus -- minimize or eliminate uses
	input lb_clk,
	input lb_strobe,
	input lb_rd,
	input [23:0] lb_addr,
	input [31:0] lb_dout,

	// clocks for frequency and phase measurement
	input U1_clkout3,
	input U2_clk_div_bufg,
	input U2_clk_div_bufr,
	input U3_clk_div_bufr,
	input bmb7_U7_clk4xout,
	input U4_dco_clk_out,

	// passed out to prc.v
	output U18_clk_in,
	output U33U1_pwr_sync,
	output [7:0] U2_idelay_ld,
	output [7:0] U3_idelay_ld,
	output [39:0] U2_idelay_value_in,
	output [39:0] U3_idelay_value_in,
	output        U15_spi_start,
	output        U15_spi_read,
	output [15:0] U15_spi_data,
	output [15:0] U15_spi_addr,
	output        U18_spi_start,
	output        U18_spi_read,
	output [23:0] U18_spi_data,
	output  [7:0] U18_spi_addr,
	output U4_reset,
	output mmcm_reset,
	input mmcm_locked,
	output U33U1_pwr_en,
	output idelayctrl_reset,

	// llspi physical I/O
	output U2_pdwn,
	output U3_pdwn,
	output U2_sclk_in,
	inout U4_sdio_inout,
	output U1_leuwire_in,
	output U27dir,
	output U2_csb_in,
	output U3_csb_in,
	output U4_csb_in,
	input U4_sdo_out,
	input U15_miso_out,
	input U18_miso_out,
	input llspi_sdi,
	output llspi_sdo,
	// slightly less physical
	output U2_clk_reset,
	output U3_clk_reset,
	output [7:0] U2_bitslip,
	output [7:0] U3_bitslip,
	output U2_iserdes_reset,
	output U3_iserdes_reset,
	output rawadc_trig_x,

	// 8 channels high-speed 16-bit parallel ADC data
	input adc_clk,
	input [127:0] adc_data,

	// outputs to host read register map
	output [31:0] banyan_status,
	output [15:0] phasex_dout,
	output [31:0] phase_status_U2,
	output [31:0] phase_status_U3,
	output  [0:0] phasex_ready,
	output  [0:0] phasex_present,
	output [7:0] llspi_status,
	output [7:0] llspi_result,
	output  [6:0] idelay_mirror_val,  // special
	output  [7:0] scanner_result_val,  // special
	output [31:0] banyan_data,  // special
	output [27:0] frequency,
	output [27:0] frequency_4xout,
	output [27:0] frequency_clkout3,
	output [27:0] frequency_dac_dco,
	output [1:0] clk_status,

	// software-settable
	input [31:0] periph_config,    // external
	input [15:0] bitslip,          // external
	input [1:0] U15_spi_read_and_start_r,  // external
	//input        U15_spi_read_r,   // external
	input [31:0] U15_spi_data_addr_r,   // external
	//input [15:0] U15_spi_addr_r,   // external
	input [1:0] U18_spi_read_and_start_r,  // external
	//input        U18_spi_read_r,   // external
	input [31:0] U18_spi_data_addr_r,   // external
	//input  [7:0] U18_spi_addr_r,   // external
	input        U2_clk_reset_r,   // external
	input        U3_clk_reset_r,   // external
	input        U2_iserdes_reset_r, // external
	input        U3_iserdes_reset_r, // external
	input        U4_reset_r,         // external
	input        mmcm_reset_r,       // external
	input        idelayctrl_reset_r, // external
	// lb_clk domain
	input [7:0] banyan_mask, // external
	input phasex_trig, // external single-cycle
	input llspi_we,  // external we-strobe
	input llspi_re,  // -- external strobe
	input clk_status_we,  // external we-strobe
	input [4:0] scanner_debug, // external
	input autoset_enable,  // -- external
	input scan_trigger,  // -- external single-cycle
	input scan_trigger_we,  // external we-strobe
	// lb_clk domain, but only because I flag_xdomain to adc_clk
	input rawadc_trig,  // external single-cycle
	// adc_clk domain
	input [9:0] sync_ad7794_cset,  // external
	input [5:0] sync_tps62210_cset  // external
);

// Propagate these (mirrored) host-settable registers to output ports of this module
assign U15_spi_start = U15_spi_read_and_start_r[0];
assign U15_spi_read = U15_spi_read_and_start_r[1];
assign U15_spi_data = U15_spi_data_addr_r[31:16];
assign U15_spi_addr = U15_spi_data_addr_r[15:0];
assign U18_spi_start = U18_spi_read_and_start_r[0];
assign U18_spi_read = U18_spi_read_and_start_r[1];
assign U18_spi_data = U18_spi_data_addr_r[31:8];
assign U18_spi_addr = U18_spi_data_addr_r[7:0];
assign U2_clk_reset = U2_clk_reset_r;
assign U3_clk_reset = U3_clk_reset_r;

assign U2_bitslip = bitslip[7:0];
assign U2_pdwn = periph_config[1];
assign U2_iserdes_reset = U2_iserdes_reset_r;
assign U3_bitslip = bitslip[15:8];
assign U3_pdwn = periph_config[1];
assign U3_iserdes_reset = U3_iserdes_reset_r;

assign U4_reset = U4_reset_r;
assign mmcm_reset = mmcm_reset_r;
assign U33U1_pwr_en = periph_config[0];
assign idelayctrl_reset = idelayctrl_reset_r;

`define CONFIG_LLSPI
`ifdef CONFIG_LLSPI
wire [8:0] host_din = lb_dout[8:0];
llspi llspi(
	.clk(lb_clk),
	// Physical FMC pins connected to digitizer board
	.P2_SCLK(U2_sclk_in),//bus_digitizer_U4[26]),
	.P2_SDI(U4_sdio_inout),//bus_digitizer_U4[0]),
	.P2_LMK_LEuWire(U1_leuwire_in),//bus_digitizer_U1[5]),
//    .P2_ADC_SDIO(U23_sdio_inout),//bus_digitizer_U4[1]),
	.sdi(llspi_sdi),
	.sdo(llspi_sdo),
	.P2_ADC_SDIO_DIR(U27dir),
	.P2_ADC_CSB_0(U2_csb_in),//bus_digitizer_U2[22]),
	.P2_ADC_CSB_1(U3_csb_in),//bus_digitizer_U3[11]),
	.P2_DAC_CSB(U4_csb_in),//bus_digitizer_U4[19]),
	.P2_DAC_SDO(U4_sdo_out),//bus_digitizer_U4[12]),
`ifdef POLL_WITH_LLSPI
// Following four llspi outputs can be left unused if
// llspi isn't driving the chips
	.P2_POLL_SCLK(U18_sclk_in),  // Y5
	.P2_POLL_MOSI(U18_mosi_in),  // V19
	.P2_AMC7823_SPI_SS(U15_ss_in),  // AB20
	.P2_AD7794_CSb(U18_ss_in),  // AE17
`endif
// OK to attach the following two llspi input pins even if
// llspi isn't driving the chips; no floating-input warnings this way
	.P2_AMC7823_SPI_MISO(U15_miso_out),//bus_digitizer_U15[1]),  // AB19
	.P2_AD7794_DOUT(U18_miso_out),//bus_digitizer_U18[1]),  // AF17
	// Host write port
	.host_din(host_din),// assign host_din = lb_dout[8:0]),
	.host_we(llspi_we),
	// Status made available to host
	.status(llspi_status),
	// Host read port
	.result_re(llspi_re),
	.host_result(llspi_result)
);
`endif

// MMCM status tracking, should detect if we ever lost clocks since setting up
// status = 0   on reset
// status = 1   set up, frozen
// status = 2   verified with PRNG
reg [1:0] clk_status_r=0;
always @(posedge lb_clk) begin
	if (clk_status_we) begin
		if (lb_dout[0]) clk_status_r <= 1;
		if (lb_dout[1] & (clk_status_r==1)) clk_status_r <= 2;
	end
	if (~mmcm_locked) clk_status_r <= 0;
end
assign clk_status = clk_status_r;

// Change clock domains for the rawadc_trig command, from lb_clk to adc_clk
flag_xdomain rawadc_trig_xdomain (.clk1(lb_clk), .flagin_clk1(rawadc_trig),
	.clk2(adc_clk), .flagout_clk2(rawadc_trig_x));

// 16 idelay registers mapped to lb_addr 112-127
// See idelay_base in static_prc_regmap.json
wire scan_running;
wire [3:0] hw_addr;
wire [4:0] hw_data;
wire hw_strobe;
wire [7:0] scanner_banyan_mask;
wire [2:0] scanner_adc_num;  // not used
wire [127:0] permuted_data;  // from banyan_mem
wire [15:0] scanner_adc_val = permuted_data[15:0];
wire lb_idelay_write = lb_strobe & ~lb_rd & (lb_addr[23:4] == 7);
idelay_scanner #(.use_decider(1)) scanner(
	.lb_clk(lb_clk), .lb_addr(lb_addr[3:0]), .lb_data(lb_dout[4:0]),
	.lb_id_write(lb_idelay_write),
	.scan_trigger(scan_trigger), .autoset_enable(autoset_enable),
	.scan_running(scan_running),
	.ro_clk(lb_clk), .ro_addr(lb_addr[10:0]),
	.mirror_val(idelay_mirror_val), .result_val(scanner_result_val),
	.debug_sel(scanner_debug[4]), .debug_addr(scanner_debug[3:0]),
	.hw_addr(hw_addr), .hw_data(hw_data), .hw_strobe(hw_strobe),
	.banyan_mask(scanner_banyan_mask), .adc_num(scanner_adc_num),
	.adc_clk(adc_clk), .adc_val(scanner_adc_val)
);

// process the output hw_ bus from idelay_scanner, sending to IDELAYE2
reg [4:0] idelay_hold=0;
reg [3:0] idelay_addr=0;
reg [1:0] idelay_sr=0;
//wire idelay_stb0 = lb_strobe & ~lb_rd &(lb_addr[23:4] == 7);
wire idelay_stb0 = hw_strobe;
// This logic is extra-fake because we don't have access to the clock used by IDELAYE2.
// Just hope we get at least one such edge every two lb_clk periods.
always @(posedge lb_clk) begin
	idelay_sr <= {idelay_sr[0],idelay_stb0};
	if (idelay_stb0) begin
		idelay_addr <= hw_addr;  //   x x A A A A x x
		idelay_hold <= hw_data;  //   x x D D D D x x
		//  idelay_stb0               __--_________
		//  idelay_stb_mask[n]        ______----_____
	end
end
reg [15:0] idelay_stb_mask=0;
genvar ixd;
generate for (ixd=0; ixd<16; ixd=ixd+1) begin: gixd
	always @(posedge lb_clk) idelay_stb_mask[ixd] <= |idelay_sr & (idelay_addr == (15-ixd));
end endgenerate
assign U2_idelay_ld = idelay_stb_mask[7:0];
assign U3_idelay_ld = idelay_stb_mask[15:8];
assign U2_idelay_value_in = {8{idelay_hold}};
assign U3_idelay_value_in = {8{idelay_hold}};

`define CONFIG_SYNC_GEN
`ifdef CONFIG_SYNC_GEN
// This is sloppy use of clock domains for sync_ad7794_cset and sync_tps62210_cset
sync_generate #(.cw(10), .minc(256)) sync_ad7794(.clk(adc_clk),
	.cset(sync_ad7794_cset), .sync(U18_clk_in));
sync_generate #(.cw(6), .minc(32)) sync_tps62210(.clk(adc_clk),
	.cset(sync_tps62210_cset), .sync(U33U1_pwr_sync));
`else
assign U18_clk_in = 0;
assign U33U1_pwr_sync = 0;
`endif

freq_count freq_count          (.clk(U3_clk_div_bufr), .usbclk(lb_clk), .frequency(frequency));
freq_count freq_count_clk4xout (.clk(bmb7_U7_clk4xout),.usbclk(lb_clk), .frequency(frequency_4xout));
freq_count freq_count_clkout3  (.clk(U1_clkout3),      .usbclk(lb_clk), .frequency(frequency_clkout3));
freq_count freq_count_dac_dco  (.clk(U4_dco_clk_out),  .usbclk(lb_clk), .frequency(frequency_dac_dco));


`define CONFIG_PHASEX
`ifdef CONFIG_PHASEX
assign phasex_present = 1;
phasex #(.aw(10)) phasex(.uclk1(U2_clk_div_bufg), .uclk2(U3_clk_div_bufr), .sclk(bmb7_U7_clk4xout),
	.rclk(lb_clk), .trig(phasex_trig), .ready(phasex_ready),
	.addr(lb_addr[9:0]), .dout(phasex_dout));
`else
assign phasex_present = 0;
assign phasex_ready = 0;
assign phasex_dout = 0;
`endif

`define CONFIG_PHASE_DIFF
`ifdef CONFIG_PHASE_DIFF
// Measure the phases of the two BUFR outputs relative to adc_clk (U2's BUFR after MMCM and BUFG)
wire [12:0] clk_phase_diff_out_U2,  clk_phase_diff_out_U3;
wire [13:0] clk_phase_diff_freq_U2, clk_phase_diff_freq_U3;
wire        clk_phase_diff_err_U2,  clk_phase_diff_err_U3;
phase_diff phase_diff_U2(.uclk1(U2_clk_div_bufg), .uclk2(U2_clk_div_bufr), .sclk(bmb7_U7_clk4xout),
	.rclk(lb_clk), .phdiff_out(clk_phase_diff_out_U2),
	.vfreq_out(clk_phase_diff_freq_U2), .err(clk_phase_diff_err_U2));
assign phase_status_U2 = {clk_phase_diff_err_U2,clk_phase_diff_freq_U2,4'b0,clk_phase_diff_out_U2};
phase_diff phase_diff_U3(.uclk1(U2_clk_div_bufg), .uclk2(U3_clk_div_bufr), .sclk(bmb7_U7_clk4xout),
	.rclk(lb_clk), .phdiff_out(clk_phase_diff_out_U3),
	.vfreq_out(clk_phase_diff_freq_U3), .err(clk_phase_diff_err_U3));
assign phase_status_U3 = {clk_phase_diff_err_U3,clk_phase_diff_freq_U3,4'b0,clk_phase_diff_out_U3};
`else
assign phase_status_U2 = 0;
assign phase_status_U3 = 0;
`endif

`define CONFIG_BANYAN
`ifdef CONFIG_BANYAN
// Banyan-routed memory, simple one-shot fill for now
parameter banyan_aw = 13;  // 8 blocks of RAM, each 8K x 16
reg banyan_run=0, banyan_run_d=0;
wire rollover, full;
wire [banyan_aw+3-1:0] pointer;
always @(posedge adc_clk) begin
	if (rawadc_trig_x | rollover) banyan_run <= rawadc_trig_x;
	banyan_run_d <= banyan_run;
end
// Control routed through idelay_scanner
reg [7:0] actual_banyan_mask=0;
always @(posedge lb_clk) actual_banyan_mask <= scan_running ? scanner_banyan_mask : banyan_mask;
// banyan_mask must be provided to banyan_mem in the adc_clk domain, otherwise the
// synthesizer will rightfully complain that timing analysis is impossible.
reg [7:0] banyan_mask_x=0;
always @(posedge adc_clk) banyan_mask_x <= actual_banyan_mask;

// Gloss over the fact that actual_banyan_mask crosses clock domains
//wire [127:0] banyan_adc = {U2DD, U2DC, U2DB, U2DA, U3DD, U3DC, U3DB, U3DA};
banyan_mem #(.aw(banyan_aw), .dw(16)) banyan_mem(.clk(adc_clk),
	.adc_data(adc_data), .banyan_mask(banyan_mask_x),
	.reset(rawadc_trig_x), .run(banyan_run),
	.pointer(pointer), .rollover(rollover), .full(full),
	.permuted_data(permuted_data),
	.ro_clk(lb_clk), .ro_addr(lb_addr[banyan_aw+3-1:0]), .ro_data(banyan_data[15:0]), .ro_data2(banyan_data[31:16])
);
// Output status can be expected to cross clock domains.
// pointer readout is only intended to be valid if ~banyan_run.
// Stretch the reported run signal to guarantee that validity rule.
wire banyan_run_s = banyan_run_d | banyan_run;
wire [5:0] banyan_aw_fix = banyan_aw;
wire [19:0] pointer_fix = pointer;
// Abuse this register a little by adding the idelay_scanner status.
// Not so bad, because that scanner depends on data provided by the banyan switch.
assign banyan_status = {banyan_run_s, full, banyan_aw_fix, 2'b0, autoset_enable, scan_running, pointer_fix};
`else
assign banyan_status = 0;
assign banyan_data = 0;
assign permuted_data = 0;
`endif

endmodule
